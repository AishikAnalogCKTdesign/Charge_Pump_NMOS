* E:\ESIM\Hackathon_Charge_Pump\Hackathon_Charge_Pump.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/02/24 01:13:09

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /

.lib "E:\ESIM\Hackathon_Charge_Pump\sky130_fd_pr\models\sky130.lib.spice" tt

XM1  Net-_XM1-Pad1_ Net-_XM1-Pad2_ Net-_C1-Pad2_ GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.50		
XM2  Net-_C1-Pad2_ Net-_XM2-Pad2_ GND GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.50		
XM3  Output_Port Net-_XM3-Pad2_ Net-_C1-Pad1_ GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.50		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 10u		
C2  Output_Port GND 1m		
v3  Net-_XM2-Pad2_ GND pulse		
v4  Net-_XM4-Pad2_ GND pulse		
v2  Net-_XM1-Pad2_ GND pulse		
v5  Net-_XM3-Pad2_ GND pulse		
V1  Net-_XM1-Pad1_ GND 5		
XM4  Net-_C1-Pad1_ Net-_XM4-Pad2_ Net-_XM1-Pad1_ GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.50		

.end
